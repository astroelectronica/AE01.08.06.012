.title KiCad schematic
.include "models/XLamp-XML-spice.txt"
V1 /IN 0 {VIN}
D1 /IN /1 XM
D2 /IN /1 XM
D3 /1 /2 XM
D4 /1 /2 XM
D5 /2 /3 XM
D6 /2 /3 XM
D7 /3 /4 XM
D8 /3 /4 XM
D9 /4 /5 XM
D10 /4 /5 XM
D11 /5 /6 XM
D12 /5 /6 XM
D13 /6 /7 XM
D14 /6 /7 XM
D15 /7 /8 XM
D16 /7 /8 XM
D17 /8 /9 XM
D18 /8 /9 XM
D19 /9 /10 XM
D20 /9 /10 XM
D21 /10 /11 XM
D22 /10 /11 XM
D23 /11 /12 XM
D24 /11 /12 XM
D25 /12 /13 XM
D26 /12 /13 XM
D27 /13 /14 XM
D28 /13 /14 XM
D29 /14 /15 XM
D30 /14 /15 XM
D31 /15 /16 XM
D32 /15 /16 XM
D33 /16 /17 XM
D34 /16 /17 XM
D35 /17 /18 XM
D36 /17 /18 XM
D37 /18 /19 XM
D38 /18 /19 XM
D39 /19 /20 XM
D40 /19 /20 XM
D41 /20 0 XM
D42 /20 0 XM
.end
